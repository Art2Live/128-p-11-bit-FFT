`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01.11.2020 21:33:43
// Design Name: 
// Module Name: FFTv2_TB
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module FFTv2_TB(

    );
    reg clk,res;
    reg   signed [10:0] In128;  // sfix11_En6
  reg   signed [10:0] In129;  // sfix11_En6
  reg   signed [10:0] In130;  // sfix11_En6
  reg   signed [10:0] In131;  // sfix11_En6
  reg   signed [10:0] In132;  // sfix11_En6
  reg   signed [10:0] In133;  // sfix11_En6
  reg   signed [10:0] In134;  // sfix11_En6
  reg   signed [10:0] In135;  // sfix11_En6
  reg   signed [10:0] In136;  // sfix11_En6
  reg   signed [10:0] In137;  // sfix11_En6
  reg   signed [10:0] In138;  // sfix11_En6
  reg   signed [10:0] In139;  // sfix11_En6
  reg   signed [10:0] In140;  // sfix11_En6
  reg   signed [10:0] In141;  // sfix11_En6
  reg   signed [10:0] In142;  // sfix11_En6
  reg   signed [10:0] In143;  // sfix11_En6
  reg   signed [10:0] In144;  // sfix11_En6
  reg   signed [10:0] In145;  // sfix11_En6
  reg   signed [10:0] In146;  // sfix11_En6
  reg   signed [10:0] In147;  // sfix11_En6
  reg   signed [10:0] In148;  // sfix11_En6
  reg   signed [10:0] In149;  // sfix11_En6
  reg   signed [10:0] In150;  // sfix11_En6
  reg   signed [10:0] In151;  // sfix11_En6
  reg   signed [10:0] In152;  // sfix11_En6
  reg   signed [10:0] In153;  // sfix11_En6
  reg   signed [10:0] In154;  // sfix11_En6
  reg   signed [10:0] In155;  // sfix11_En6
  reg   signed [10:0] In156;  // sfix11_En6
  reg   signed [10:0] In157;  // sfix11_En6
  reg   signed [10:0] In158;  // sfix11_En6
  reg   signed [10:0] In159;  // sfix11_En6
  reg   signed [10:0] In160;  // sfix11_En6
  reg   signed [10:0] In161;  // sfix11_En6
  reg   signed [10:0] In162;  // sfix11_En6
  reg   signed [10:0] In163;  // sfix11_En6
  reg   signed [10:0] In164;  // sfix11_En6
  reg   signed [10:0] In165;  // sfix11_En6
  reg   signed [10:0] In166;  // sfix11_En6
  reg   signed [10:0] In167;  // sfix11_En6
  reg   signed [10:0] In168;  // sfix11_En6
  reg   signed [10:0] In169;  // sfix11_En6
  reg   signed [10:0] In170;  // sfix11_En6
  reg   signed [10:0] In171;  // sfix11_En6
  reg   signed [10:0] In172;  // sfix11_En6
  reg   signed [10:0] In173;  // sfix11_En6
  reg   signed [10:0] In174;  // sfix11_En6
  reg   signed [10:0] In175;  // sfix11_En6
  reg   signed [10:0] In176;  // sfix11_En6
  reg   signed [10:0] In177;  // sfix11_En6
  reg   signed [10:0] In178;  // sfix11_En6
  reg   signed [10:0] In179;  // sfix11_En6
  reg   signed [10:0] In180;  // sfix11_En6
  reg   signed [10:0] In181;  // sfix11_En6
  reg   signed [10:0] In182;  // sfix11_En6
  reg   signed [10:0] In183;  // sfix11_En6
  reg   signed [10:0] In184;  // sfix11_En6
  reg   signed [10:0] In185;  // sfix11_En6
  reg   signed [10:0] In186;  // sfix11_En6
  reg   signed [10:0] In187;  // sfix11_En6
  reg   signed [10:0] In188;  // sfix11_En6
  reg   signed [10:0] In189;  // sfix11_En6
  reg   signed [10:0] In190;  // sfix11_En6
  reg   signed [10:0] In191;  // sfix11_En6
  reg   signed [10:0] In192;  // sfix11_En6
  reg   signed [10:0] In193;  // sfix11_En6
  reg   signed [10:0] In194;  // sfix11_En6
  reg   signed [10:0] In195;  // sfix11_En6
  reg   signed [10:0] In196;  // sfix11_En6
  reg   signed [10:0] In197;  // sfix11_En6
  reg   signed [10:0] In198;  // sfix11_En6
  reg   signed [10:0] In199;  // sfix11_En6
  reg   signed [10:0] In200;  // sfix11_En6
  reg   signed [10:0] In201;  // sfix11_En6
  reg   signed [10:0] In202;  // sfix11_En6
  reg   signed [10:0] In203;  // sfix11_En6
  reg   signed [10:0] In204;  // sfix11_En6
  reg   signed [10:0] In205;  // sfix11_En6
  reg   signed [10:0] In206;  // sfix11_En6
  reg   signed [10:0] In207;  // sfix11_En6
  reg   signed [10:0] In208;  // sfix11_En6
  reg   signed [10:0] In209;  // sfix11_En6
  reg   signed [10:0] In210;  // sfix11_En6
  reg   signed [10:0] In211;  // sfix11_En6
  reg   signed [10:0] In212;  // sfix11_En6
  reg   signed [10:0] In213;  // sfix11_En6
  reg   signed [10:0] In214;  // sfix11_En6
  reg   signed [10:0] In215;  // sfix11_En6
  reg   signed [10:0] In216;  // sfix11_En6
  reg   signed [10:0] In217;  // sfix11_En6
  reg   signed [10:0] In218;  // sfix11_En6
  reg   signed [10:0] In219;  // sfix11_En6
  reg   signed [10:0] In220;  // sfix11_En6
  reg   signed [10:0] In221;  // sfix11_En6
  reg   signed [10:0] In222;  // sfix11_En6
  reg   signed [10:0] In223;  // sfix11_En6
  reg   signed [10:0] In224;  // sfix11_En6
  reg   signed [10:0] In225;  // sfix11_En6
  reg   signed [10:0] In226;  // sfix11_En6
  reg   signed [10:0] In227;  // sfix11_En6
  reg   signed [10:0] In228;  // sfix11_En6
  reg   signed [10:0] In229;  // sfix11_En6
  reg   signed [10:0] In230;  // sfix11_En6
  reg   signed [10:0] In231;  // sfix11_En6
  reg   signed [10:0] In232;  // sfix11_En6
  reg   signed [10:0] In233;  // sfix11_En6
  reg   signed [10:0] In234;  // sfix11_En6
  reg   signed [10:0] In235;  // sfix11_En6
  reg   signed [10:0] In236;  // sfix11_En6
  reg   signed [10:0] In237;  // sfix11_En6
  reg   signed [10:0] In238;  // sfix11_En6
  reg   signed [10:0] In239;  // sfix11_En6
  reg   signed [10:0] In240;  // sfix11_En6
  reg   signed [10:0] In241;  // sfix11_En6
  reg   signed [10:0] In242;  // sfix11_En6
  reg   signed [10:0] In243;  // sfix11_En6
  reg   signed [10:0] In244;  // sfix11_En6
  reg   signed [10:0] In245;  // sfix11_En6
  reg   signed [10:0] In246;  // sfix11_En6
  reg   signed [10:0] In247;  // sfix11_En6
  reg   signed [10:0] In248;  // sfix11_En6
  reg   signed [10:0] In249;  // sfix11_En6
  reg   signed [10:0] In250;  // sfix11_En6
  reg   signed [10:0] In251;  // sfix11_En6
  reg   signed [10:0] In252;  // sfix11_En6
  reg   signed [10:0] In253;  // sfix11_En6
  reg   signed [10:0] In254;  // sfix11_En6
  reg   signed [10:0] In255;  // sfix11_En6
wire  signed [10:0] Out1_re;  // sfix11
  wire  signed [10:0] Out1_im;  // sfix11
  wire  signed [10:0] Out2_re;  // sfix11
  wire  signed [10:0] Out2_im;  // sfix11
  wire  signed [10:0] Out3_re;  // sfix11
  wire  signed [10:0] Out3_im;  // sfix11
  wire  signed [10:0] Out4_re;  // sfix11
  wire  signed [10:0] Out4_im;  // sfix11
  wire  signed [10:0] Out5_re;  // sfix11
  wire  signed [10:0] Out5_im;  // sfix11
  wire  signed [10:0] Out6_re;  // sfix11
  wire  signed [10:0] Out6_im;  // sfix11
  wire  signed [10:0] Out7_re;  // sfix11
  wire  signed [10:0] Out7_im;  // sfix11
  wire  signed [10:0] Out8_re;  // sfix11
  wire  signed [10:0] Out8_im;  // sfix11
  wire  signed [10:0] Out9_re;  // sfix11
  wire  signed [10:0] Out9_im;  // sfix11
  wire  signed [10:0] Out10_re;  // sfix11
  wire  signed [10:0] Out10_im;  // sfix11
  wire  signed [10:0] Out11_re;  // sfix11
  wire  signed [10:0] Out11_im;  // sfix11
  wire  signed [10:0] Out12_re;  // sfix11
  wire  signed [10:0] Out12_im;  // sfix11
  wire  signed [10:0] Out13_re;  // sfix11
  wire  signed [10:0] Out13_im;  // sfix11
  wire  signed [10:0] Out14_re;  // sfix11
  wire  signed [10:0] Out14_im;  // sfix11
  wire  signed [10:0] Out15_re;  // sfix11
  wire  signed [10:0] Out15_im;  // sfix11
  wire  signed [10:0] Out16_re;  // sfix11
  wire  signed [10:0] Out16_im;  // sfix11
  wire  signed [10:0] Out17_re;  // sfix11
  wire  signed [10:0] Out17_im;  // sfix11
  wire  signed [10:0] Out18_re;  // sfix11
  wire  signed [10:0] Out18_im;  // sfix11
  wire  signed [10:0] Out19_re;  // sfix11
  wire  signed [10:0] Out19_im;  // sfix11
  wire  signed [10:0] Out20_re;  // sfix11
  wire  signed [10:0] Out20_im;  // sfix11
  wire  signed [10:0] Out21_re;  // sfix11
  wire  signed [10:0] Out21_im;  // sfix11
  wire  signed [10:0] Out22_re;  // sfix11
  wire  signed [10:0] Out22_im;  // sfix11
  wire  signed [10:0] Out23_re;  // sfix11
  wire  signed [10:0] Out23_im;  // sfix11
  wire  signed [10:0] Out24_re;  // sfix11
  wire  signed [10:0] Out24_im;  // sfix11
  wire  signed [10:0] Out25_re;  // sfix11
  wire  signed [10:0] Out25_im;  // sfix11
  wire  signed [10:0] Out26_re;  // sfix11
  wire  signed [10:0] Out26_im;  // sfix11
  wire  signed [10:0] Out27_re;  // sfix11
  wire  signed [10:0] Out27_im;  // sfix11
  wire  signed [10:0] Out28_re;  // sfix11
  wire  signed [10:0] Out28_im;  // sfix11
  wire  signed [10:0] Out29_re;  // sfix11
  wire  signed [10:0] Out29_im;  // sfix11
  wire  signed [10:0] Out30_re;  // sfix11
  wire  signed [10:0] Out30_im;  // sfix11
  wire  signed [10:0] Out31_re;  // sfix11
  wire  signed [10:0] Out31_im;  // sfix11
  wire  signed [10:0] Out32_re;  // sfix11
  wire  signed [10:0] Out32_im;  // sfix11
  wire  signed [10:0] Out33_re;  // sfix11
  wire  signed [10:0] Out33_im;  // sfix11
  wire  signed [10:0] Out34_re;  // sfix11
  wire  signed [10:0] Out34_im;  // sfix11
  wire  signed [10:0] Out35_re;  // sfix11
  wire  signed [10:0] Out35_im;  // sfix11
  wire  signed [10:0] Out36_re;  // sfix11
  wire  signed [10:0] Out36_im;  // sfix11
  wire  signed [10:0] Out37_re;  // sfix11
  wire  signed [10:0] Out37_im;  // sfix11
  wire  signed [10:0] Out38_re;  // sfix11
  wire  signed [10:0] Out38_im;  // sfix11
  wire  signed [10:0] Out39_re;  // sfix11
  wire  signed [10:0] Out39_im;  // sfix11
  wire  signed [10:0] Out40_re;  // sfix11
  wire  signed [10:0] Out40_im;  // sfix11
  wire  signed [10:0] Out41_re;  // sfix11
  wire  signed [10:0] Out41_im;  // sfix11
  wire  signed [10:0] Out42_re;  // sfix11
  wire  signed [10:0] Out42_im;  // sfix11
  wire  signed [10:0] Out43_re;  // sfix11
  wire  signed [10:0] Out43_im;  // sfix11
  wire  signed [10:0] Out44_re;  // sfix11
  wire  signed [10:0] Out44_im;  // sfix11
  wire  signed [10:0] Out45_re;  // sfix11
  wire  signed [10:0] Out45_im;  // sfix11
  wire  signed [10:0] Out46_re;  // sfix11
  wire  signed [10:0] Out46_im;  // sfix11
  wire  signed [10:0] Out47_re;  // sfix11
  wire  signed [10:0] Out47_im;  // sfix11
  wire  signed [10:0] Out48_re;  // sfix11
  wire  signed [10:0] Out48_im;  // sfix11
  wire  signed [10:0] Out49_re;  // sfix11
  wire  signed [10:0] Out49_im;  // sfix11
  wire  signed [10:0] Out50_re;  // sfix11
  wire  signed [10:0] Out50_im;  // sfix11
  wire  signed [10:0] Out51_re;  // sfix11
  wire  signed [10:0] Out51_im;  // sfix11
  wire  signed [10:0] Out52_re;  // sfix11
  wire  signed [10:0] Out52_im;  // sfix11
  wire  signed [10:0] Out53_re;  // sfix11
  wire  signed [10:0] Out53_im;  // sfix11
  wire  signed [10:0] Out54_re;  // sfix11
  wire  signed [10:0] Out54_im;  // sfix11
  wire  signed [10:0] Out55_re;  // sfix11
  wire  signed [10:0] Out55_im;  // sfix11
  wire  signed [10:0] Out56_re;  // sfix11
  wire  signed [10:0] Out56_im;  // sfix11
  wire  signed [10:0] Out57_re;  // sfix11
  wire  signed [10:0] Out57_im;  // sfix11
  wire  signed [10:0] Out58_re;  // sfix11
  wire  signed [10:0] Out58_im;  // sfix11
  wire  signed [10:0] Out59_re;  // sfix11
  wire  signed [10:0] Out59_im;  // sfix11
  wire  signed [10:0] Out60_re;  // sfix11
  wire  signed [10:0] Out60_im;  // sfix11
  wire  signed [10:0] Out61_re;  // sfix11
  wire  signed [10:0] Out61_im;  // sfix11
  wire  signed [10:0] Out62_re;  // sfix11
  wire  signed [10:0] Out62_im;  // sfix11
  wire  signed [10:0] Out63_re;  // sfix11
  wire  signed [10:0] Out63_im;  // sfix11
  wire  signed [10:0] Out64_re;  // sfix11
  wire  signed [10:0] Out64_im;  // sfix11
  wire  signed [10:0] Out65_re;  // sfix11
  wire  signed [10:0] Out65_im;  // sfix11
  wire  signed [10:0] Out66_re;  // sfix11
  wire  signed [10:0] Out66_im;  // sfix11
  wire  signed [10:0] Out67_re;  // sfix11
  wire  signed [10:0] Out67_im;  // sfix11
  wire  signed [10:0] Out68_re;  // sfix11
  wire  signed [10:0] Out68_im;  // sfix11
  wire  signed [10:0] Out69_re;  // sfix11
  wire  signed [10:0] Out69_im;  // sfix11
  wire  signed [10:0] Out70_re;  // sfix11
  wire  signed [10:0] Out70_im;  // sfix11
  wire  signed [10:0] Out71_re;  // sfix11
  wire  signed [10:0] Out71_im;  // sfix11
  wire  signed [10:0] Out72_re;  // sfix11
  wire  signed [10:0] Out72_im;  // sfix11
  wire  signed [10:0] Out73_re;  // sfix11
  wire  signed [10:0] Out73_im;  // sfix11
  wire  signed [10:0] Out74_re;  // sfix11
  wire  signed [10:0] Out74_im;  // sfix11
  wire  signed [10:0] Out75_re;  // sfix11
  wire  signed [10:0] Out75_im;  // sfix11
  wire  signed [10:0] Out76_re;  // sfix11
  wire  signed [10:0] Out76_im;  // sfix11
  wire  signed [10:0] Out77_re;  // sfix11
  wire  signed [10:0] Out77_im;  // sfix11
  wire  signed [10:0] Out78_re;  // sfix11
  wire  signed [10:0] Out78_im;  // sfix11
  wire  signed [10:0] Out79_re;  // sfix11
  wire  signed [10:0] Out79_im;  // sfix11
  wire  signed [10:0] Out80_re;  // sfix11
  wire  signed [10:0] Out80_im;  // sfix11
  wire  signed [10:0] Out81_re;  // sfix11
  wire  signed [10:0] Out81_im;  // sfix11
  wire  signed [10:0] Out82_re;  // sfix11
  wire  signed [10:0] Out82_im;  // sfix11
  wire  signed [10:0] Out83_re;  // sfix11
  wire  signed [10:0] Out83_im;  // sfix11
  wire  signed [10:0] Out84_re;  // sfix11
  wire  signed [10:0] Out84_im;  // sfix11
  wire  signed [10:0] Out85_re;  // sfix11
  wire  signed [10:0] Out85_im;  // sfix11
  wire  signed [10:0] Out86_re;  // sfix11
  wire  signed [10:0] Out86_im;  // sfix11
  wire  signed [10:0] Out87_re;  // sfix11
  wire  signed [10:0] Out87_im;  // sfix11
  wire  signed [10:0] Out88_re;  // sfix11
  wire  signed [10:0] Out88_im;  // sfix11
  wire  signed [10:0] Out89_re;  // sfix11
  wire  signed [10:0] Out89_im;  // sfix11
  wire  signed [10:0] Out90_re;  // sfix11
  wire  signed [10:0] Out90_im;  // sfix11
  wire  signed [10:0] Out91_re;  // sfix11
  wire  signed [10:0] Out91_im;  // sfix11
  wire  signed [10:0] Out92_re;  // sfix11
  wire  signed [10:0] Out92_im;  // sfix11
  wire  signed [10:0] Out93_re;  // sfix11
  wire  signed [10:0] Out93_im;  // sfix11
  wire  signed [10:0] Out94_re;  // sfix11
  wire  signed [10:0] Out94_im;  // sfix11
  wire  signed [10:0] Out95_re;  // sfix11
  wire  signed [10:0] Out95_im;  // sfix11
  wire  signed [10:0] Out96_re;  // sfix11
  wire  signed [10:0] Out96_im;  // sfix11
  wire  signed [10:0] Out97_re;  // sfix11
  wire  signed [10:0] Out97_im;  // sfix11
  wire  signed [10:0] Out98_re;  // sfix11
  wire  signed [10:0] Out98_im;  // sfix11
  wire  signed [10:0] Out99_re;  // sfix11
  wire  signed [10:0] Out99_im;  // sfix11
  wire  signed [10:0] Out100_re;  // sfix11
  wire  signed [10:0] Out100_im;  // sfix11
  wire  signed [10:0] Out101_re;  // sfix11
  wire  signed [10:0] Out101_im;  // sfix11
  wire  signed [10:0] Out102_re;  // sfix11
  wire  signed [10:0] Out102_im;  // sfix11
  wire  signed [10:0] Out103_re;  // sfix11
  wire  signed [10:0] Out103_im;  // sfix11
  wire  signed [10:0] Out104_re;  // sfix11
  wire  signed [10:0] Out104_im;  // sfix11
  wire  signed [10:0] Out105_re;  // sfix11
  wire  signed [10:0] Out105_im;  // sfix11
  wire  signed [10:0] Out106_re;  // sfix11
  wire  signed [10:0] Out106_im;  // sfix11
  wire  signed [10:0] Out107_re;  // sfix11
  wire  signed [10:0] Out107_im;  // sfix11
  wire  signed [10:0] Out108_re;  // sfix11
  wire  signed [10:0] Out108_im;  // sfix11
  wire  signed [10:0] Out109_re;  // sfix11
  wire  signed [10:0] Out109_im;  // sfix11
  wire  signed [10:0] Out110_re;  // sfix11
  wire  signed [10:0] Out110_im;  // sfix11
  wire  signed [10:0] Out111_re;  // sfix11
  wire  signed [10:0] Out111_im;  // sfix11
  wire  signed [10:0] Out112_re;  // sfix11
  wire  signed [10:0] Out112_im;  // sfix11
  wire  signed [10:0] Out113_re;  // sfix11
  wire  signed [10:0] Out113_im;  // sfix11
  wire  signed [10:0] Out114_re;  // sfix11
  wire  signed [10:0] Out114_im;  // sfix11
  wire  signed [10:0] Out115_re;  // sfix11
  wire  signed [10:0] Out115_im;  // sfix11
  wire  signed [10:0] Out116_re;  // sfix11
  wire  signed [10:0] Out116_im;  // sfix11
  wire  signed [10:0] Out117_re;  // sfix11
  wire  signed [10:0] Out117_im;  // sfix11
  wire  signed [10:0] Out118_re;  // sfix11
  wire  signed [10:0] Out118_im;  // sfix11
  wire  signed [10:0] Out119_re;  // sfix11
  wire  signed [10:0] Out119_im;  // sfix11
  wire  signed [10:0] Out120_re;  // sfix11
  wire  signed [10:0] Out120_im;  // sfix11
  wire  signed [10:0] Out121_re;  // sfix11
  wire  signed [10:0] Out121_im;  // sfix11
  wire  signed [10:0] Out122_re;  // sfix11
  wire  signed [10:0] Out122_im;  // sfix11
  wire  signed [10:0] Out123_re;  // sfix11
  wire  signed [10:0] Out123_im;  // sfix11
  wire  signed [10:0] Out124_re;  // sfix11
  wire  signed [10:0] Out124_im;  // sfix11
  wire  signed [10:0] Out125_re;  // sfix11
  wire  signed [10:0] Out125_im;  // sfix11
  wire  signed [10:0] Out126_re;  // sfix11
  wire  signed [10:0] Out126_im;  // sfix11
  wire  signed [10:0] Out127_re;  // sfix11
  wire  signed [10:0] Out127_im;  // sfix11
  wire  signed [10:0] Out128_re;  // sfix11
  wire  signed [10:0] Out128_im;  // sfix11 
    FFTv2 uut (  .clk(clk), .reset(res),  
    .In1(In128),  // sfix11_En6
                                          .In2(In129),  // sfix11_En6
                                          .In3(In130),  // sfix11_En6
                                          .In4(In131),  // sfix11_En6
                                          .In5(In132),  // sfix11_En6
                                          .In6(In133),  // sfix11_En6
                                          .In7(In134),  // sfix11_En6
                                          .In8(In135),  // sfix11_En6
                                          .In9(In136),  // sfix11_En6
                                          .In10(In137),  // sfix11_En6
                                          .In11(In138),  // sfix11_En6
                                          .In12(In139),  // sfix11_En6
                                          .In13(In140),  // sfix11_En6
                                          .In14(In141),  // sfix11_En6
                                          .In15(In142),  // sfix11_En6
                                          .In16(In143),  // sfix11_En6
                                          .In17(In144),  // sfix11_En6
                                          .In18(In145),  // sfix11_En6
                                          .In19(In146),  // sfix11_En6
                                          .In20(In147),  // sfix11_En6
                                          .In21(In148),  // sfix11_En6
                                          .In22(In149),  // sfix11_En6
                                          .In23(In150),  // sfix11_En6
                                          .In24(In151),  // sfix11_En6
                                          .In25(In152),  // sfix11_En6
                                          .In26(In153),  // sfix11_En6
                                          .In27(In154),  // sfix11_En6
                                          .In28(In155),  // sfix11_En6
                                          .In29(In156),  // sfix11_En6
                                          .In30(In157),  // sfix11_En6
                                          .In31(In158),  // sfix11_En6
                                          .In32(In159),  // sfix11_En6
                                          .In33(In160),  // sfix11_En6
                                          .In34(In161),  // sfix11_En6
                                          .In35(In162),  // sfix11_En6
                                          .In36(In163),  // sfix11_En6
                                          .In37(In164),  // sfix11_En6
                                          .In38(In165),  // sfix11_En6
                                          .In39(In166),  // sfix11_En6
                                          .In40(In167),  // sfix11_En6
                                          .In41(In168),  // sfix11_En6
                                          .In42(In169),  // sfix11_En6
                                          .In43(In170),  // sfix11_En6
                                          .In44(In171),  // sfix11_En6
                                          .In45(In172),  // sfix11_En6
                                          .In46(In173),  // sfix11_En6
                                          .In47(In174),  // sfix11_En6
                                          .In48(In175),  // sfix11_En6
                                          .In49(In176),  // sfix11_En6
                                          .In50(In177),  // sfix11_En6
                                          .In51(In178),  // sfix11_En6
                                          .In52(In179),  // sfix11_En6
                                          .In53(In180),  // sfix11_En6
                                          .In54(In181),  // sfix11_En6
                                          .In55(In182),  // sfix11_En6
                                          .In56(In183),  // sfix11_En6
                                          .In57(In184),  // sfix11_En6
                                          .In58(In185),  // sfix11_En6
                                          .In59(In186),  // sfix11_En6
                                          .In60(In187),  // sfix11_En6
                                          .In61(In188),  // sfix11_En6
                                          .In62(In189),  // sfix11_En6
                                          .In63(In190),  // sfix11_En6
                                          .In64(In191),  // sfix11_En6
                                          .In65(In192),  // sfix11_En6
                                          .In66(In193),  // sfix11_En6
                                          .In67(In194),  // sfix11_En6
                                          .In68(In195),  // sfix11_En6
                                          .In69(In196),  // sfix11_En6
                                          .In70(In197),  // sfix11_En6
                                          .In71(In198),  // sfix11_En6
                                          .In72(In199),  // sfix11_En6
                                          .In73(In200),  // sfix11_En6
                                          .In74(In201),  // sfix11_En6
                                          .In75(In202),  // sfix11_En6
                                          .In76(In203),  // sfix11_En6
                                          .In77(In204),  // sfix11_En6
                                          .In78(In205),  // sfix11_En6
                                          .In79(In206),  // sfix11_En6
                                          .In80(In207),  // sfix11_En6
                                          .In81(In208),  // sfix11_En6
                                          .In82(In209),  // sfix11_En6
                                          .In83(In210),  // sfix11_En6
                                          .In84(In211),  // sfix11_En6
                                          .In85(In212),  // sfix11_En6
                                          .In86(In213),  // sfix11_En6
                                          .In87(In214),  // sfix11_En6
                                          .In88(In215),  // sfix11_En6
                                          .In89(In216),  // sfix11_En6
                                          .In90(In217),  // sfix11_En6
                                          .In91(In218),  // sfix11_En6
                                          .In92(In219),  // sfix11_En6
                                          .In93(In220),  // sfix11_En6
                                          .In94(In221),  // sfix11_En6
                                          .In95(In222),  // sfix11_En6
                                          .In96(In223),  // sfix11_En6
                                          .In97(In224),  // sfix11_En6
                                          .In98(In225),  // sfix11_En6
                                          .In99(In226),  // sfix11_En6
                                          .In100(In227),  // sfix11_En6
                                          .In101(In228),  // sfix11_En6
                                          .In102(In229),  // sfix11_En6
                                          .In103(In230),  // sfix11_En6
                                          .In104(In231),  // sfix11_En6
                                          .In105(In232),  // sfix11_En6
                                          .In106(In233),  // sfix11_En6
                                          .In107(In234),  // sfix11_En6
                                          .In108(In235),  // sfix11_En6
                                          .In109(In236),  // sfix11_En6
                                          .In110(In237),  // sfix11_En6
                                          .In111(In238),  // sfix11_En6
                                          .In112(In239),  // sfix11_En6
                                          .In113(In240),  // sfix11_En6
                                          .In114(In241),  // sfix11_En6
                                          .In115(In242),  // sfix11_En6
                                          .In116(In243),  // sfix11_En6
                                          .In117(In244),  // sfix11_En6
                                          .In118(In245),  // sfix11_En6
                                          .In119(In246),  // sfix11_En6
                                          .In120(In247),  // sfix11_En6
                                          .In121(In248),  // sfix11_En6
                                          .In122(In249),  // sfix11_En6
                                          .In123(In250),  // sfix11_En6
                                          .In124(In251),  // sfix11_En6
                                          .In125(In252),  // sfix11_En6
                                          .In126(In253),  // sfix11_En6
                                          .In127(In254),  // sfix11_En6
                                          .In128(In255),  // sfix11_En6   
                                          .Out1_re(Out1_re),  
                             .Out1_im(Out1_im),  
                             .Out2_re(Out2_re),  
                             .Out2_im(Out2_im),  
                             .Out3_re(Out3_re),  
                             .Out3_im(Out3_im),  
                             .Out4_re(Out4_re),  
                             .Out4_im(Out4_im),  
                             .Out5_re(Out5_re),  
                             .Out5_im(Out5_im),  
                             .Out6_re(Out6_re),  
                             .Out6_im(Out6_im),  
                             .Out7_re(Out7_re),  
                             .Out7_im(Out7_im),  
                             .Out8_re(Out8_re),  
                             .Out8_im(Out8_im),  
                             .Out9_re(Out9_re),  
                             .Out9_im(Out9_im),  
                             .Out10_re(Out10_re),  
                             .Out10_im(Out10_im),  
                             .Out11_re(Out11_re),  
                             .Out11_im(Out11_im),  
                             .Out12_re(Out12_re),  
                             .Out12_im(Out12_im),  
                             .Out13_re(Out13_re),  
                             .Out13_im(Out13_im),  
                             .Out14_re(Out14_re),  
                             .Out14_im(Out14_im),  
                             .Out15_re(Out15_re),  
                             .Out15_im(Out15_im),  
                             .Out16_re(Out16_re),  
                             .Out16_im(Out16_im),  
                             .Out17_re(Out17_re),  
                             .Out17_im(Out17_im),  
                             .Out18_re(Out18_re),  
                             .Out18_im(Out18_im),  
                             .Out19_re(Out19_re),  
                             .Out19_im(Out19_im),  
                             .Out20_re(Out20_re),  
                             .Out20_im(Out20_im),  
                             .Out21_re(Out21_re),  
                             .Out21_im(Out21_im),  
                             .Out22_re(Out22_re),  
                             .Out22_im(Out22_im),  
                             .Out23_re(Out23_re),  
                             .Out23_im(Out23_im),  
                             .Out24_re(Out24_re),  
                             .Out24_im(Out24_im),  
                             .Out25_re(Out25_re),  
                             .Out25_im(Out25_im),  
                             .Out26_re(Out26_re),  
                             .Out26_im(Out26_im),  
                             .Out27_re(Out27_re),  
                             .Out27_im(Out27_im),  
                             .Out28_re(Out28_re),  
                             .Out28_im(Out28_im),  
                             .Out29_re(Out29_re),  
                             .Out29_im(Out29_im),  
                             .Out30_re(Out30_re),  
                             .Out30_im(Out30_im),  
                             .Out31_re(Out31_re),  
                             .Out31_im(Out31_im),  
                             .Out32_re(Out32_re),  
                             .Out32_im(Out32_im),  
                             .Out33_re(Out33_re),  
                             .Out33_im(Out33_im),  
                             .Out34_re(Out34_re),  
                             .Out34_im(Out34_im),  
                             .Out35_re(Out35_re),  
                             .Out35_im(Out35_im),  
                             .Out36_re(Out36_re),  
                             .Out36_im(Out36_im),  
                             .Out37_re(Out37_re),  
                             .Out37_im(Out37_im),  
                             .Out38_re(Out38_re),  
                             .Out38_im(Out38_im),  
                             .Out39_re(Out39_re),  
                             .Out39_im(Out39_im),  
                             .Out40_re(Out40_re),  
                             .Out40_im(Out40_im),  
                             .Out41_re(Out41_re),  
                             .Out41_im(Out41_im),  
                             .Out42_re(Out42_re),  
                             .Out42_im(Out42_im),  
                             .Out43_re(Out43_re),  
                             .Out43_im(Out43_im),  
                             .Out44_re(Out44_re),  
                             .Out44_im(Out44_im),  
                             .Out45_re(Out45_re),  
                             .Out45_im(Out45_im),  
                             .Out46_re(Out46_re),  
                             .Out46_im(Out46_im),  
                             .Out47_re(Out47_re),  
                             .Out47_im(Out47_im),  
                             .Out48_re(Out48_re),  
                             .Out48_im(Out48_im),  
                             .Out49_re(Out49_re),  
                             .Out49_im(Out49_im),  
                             .Out50_re(Out50_re),  
                             .Out50_im(Out50_im),  
                             .Out51_re(Out51_re),  
                             .Out51_im(Out51_im),  
                             .Out52_re(Out52_re),  
                             .Out52_im(Out52_im),  
                             .Out53_re(Out53_re),  
                             .Out53_im(Out53_im),  
                             .Out54_re(Out54_re),  
                             .Out54_im(Out54_im),  
                             .Out55_re(Out55_re),  
                             .Out55_im(Out55_im),  
                             .Out56_re(Out56_re),  
                             .Out56_im(Out56_im),  
                             .Out57_re(Out57_re),  
                             .Out57_im(Out57_im),  
                             .Out58_re(Out58_re),  
                             .Out58_im(Out58_im),  
                             .Out59_re(Out59_re),  
                             .Out59_im(Out59_im),  
                             .Out60_re(Out60_re),  
                             .Out60_im(Out60_im),  
                             .Out61_re(Out61_re),  
                             .Out61_im(Out61_im),  
                             .Out62_re(Out62_re),  
                             .Out62_im(Out62_im),  
                             .Out63_re(Out63_re),  
                             .Out63_im(Out63_im),  
                             .Out64_re(Out64_re),  
                             .Out64_im(Out64_im),  
                             .Out65_re(Out65_re),  
                             .Out65_im(Out65_im),  
                             .Out66_re(Out66_re),  
                             .Out66_im(Out66_im),  
                             .Out67_re(Out67_re),  
                             .Out67_im(Out67_im),  
                             .Out68_re(Out68_re),  
                             .Out68_im(Out68_im),  
                             .Out69_re(Out69_re),  
                             .Out69_im(Out69_im),  
                             .Out70_re(Out70_re),  
                             .Out70_im(Out70_im),  
                             .Out71_re(Out71_re),  
                             .Out71_im(Out71_im),  
                             .Out72_re(Out72_re),  
                             .Out72_im(Out72_im),  
                             .Out73_re(Out73_re),  
                             .Out73_im(Out73_im),  
                             .Out74_re(Out74_re),  
                             .Out74_im(Out74_im),  
                             .Out75_re(Out75_re),  
                             .Out75_im(Out75_im),  
                             .Out76_re(Out76_re),  
                             .Out76_im(Out76_im),  
                             .Out77_re(Out77_re),  
                             .Out77_im(Out77_im),  
                             .Out78_re(Out78_re),  
                             .Out78_im(Out78_im),  
                             .Out79_re(Out79_re),  
                             .Out79_im(Out79_im),  
                             .Out80_re(Out80_re),  
                             .Out80_im(Out80_im),  
                             .Out81_re(Out81_re),  
                             .Out81_im(Out81_im),  
                             .Out82_re(Out82_re),  
                             .Out82_im(Out82_im),  
                             .Out83_re(Out83_re),  
                             .Out83_im(Out83_im),  
                             .Out84_re(Out84_re),  
                             .Out84_im(Out84_im),  
                             .Out85_re(Out85_re),  
                             .Out85_im(Out85_im),  
                             .Out86_re(Out86_re),  
                             .Out86_im(Out86_im),  
                             .Out87_re(Out87_re),  
                             .Out87_im(Out87_im),  
                             .Out88_re(Out88_re),  
                             .Out88_im(Out88_im),  
                             .Out89_re(Out89_re),  
                             .Out89_im(Out89_im),  
                             .Out90_re(Out90_re),  
                             .Out90_im(Out90_im),  
                             .Out91_re(Out91_re),  
                             .Out91_im(Out91_im),  
                             .Out92_re(Out92_re),  
                             .Out92_im(Out92_im),  
                             .Out93_re(Out93_re),  
                             .Out93_im(Out93_im),  
                             .Out94_re(Out94_re),  
                             .Out94_im(Out94_im),  
                             .Out95_re(Out95_re),  
                             .Out95_im(Out95_im),  
                             .Out96_re(Out96_re),  
                             .Out96_im(Out96_im),  
                             .Out97_re(Out97_re),  
                             .Out97_im(Out97_im),  
                             .Out98_re(Out98_re),  
                             .Out98_im(Out98_im),  
                             .Out99_re(Out99_re),  
                             .Out99_im(Out99_im),  
                             .Out100_re(Out100_re),  
                             .Out100_im(Out100_im),  
                             .Out101_re(Out101_re),  
                             .Out101_im(Out101_im),  
                             .Out102_re(Out102_re),  
                             .Out102_im(Out102_im),  
                             .Out103_re(Out103_re),  
                             .Out103_im(Out103_im),  
                             .Out104_re(Out104_re),  
                             .Out104_im(Out104_im),  
                             .Out105_re(Out105_re),  
                             .Out105_im(Out105_im),  
                             .Out106_re(Out106_re),  
                             .Out106_im(Out106_im),  
                             .Out107_re(Out107_re),  
                             .Out107_im(Out107_im),  
                             .Out108_re(Out108_re),  
                             .Out108_im(Out108_im),  
                             .Out109_re(Out109_re),  
                             .Out109_im(Out109_im),  
                             .Out110_re(Out110_re),  
                             .Out110_im(Out110_im),  
                             .Out111_re(Out111_re),  
                             .Out111_im(Out111_im),  
                             .Out112_re(Out112_re),  
                             .Out112_im(Out112_im),  
                             .Out113_re(Out113_re),  
                             .Out113_im(Out113_im),  
                             .Out114_re(Out114_re),  
                             .Out114_im(Out114_im),  
                             .Out115_re(Out115_re),  
                             .Out115_im(Out115_im),  
                             .Out116_re(Out116_re),  
                             .Out116_im(Out116_im),  
                             .Out117_re(Out117_re),  
                             .Out117_im(Out117_im),  
                             .Out118_re(Out118_re),  
                             .Out118_im(Out118_im),  
                             .Out119_re(Out119_re),  
                             .Out119_im(Out119_im),  
                             .Out120_re(Out120_re),  
                             .Out120_im(Out120_im),  
                             .Out121_re(Out121_re),  
                             .Out121_im(Out121_im),  
                             .Out122_re(Out122_re),  
                             .Out122_im(Out122_im),  
                             .Out123_re(Out123_re),  
                             .Out123_im(Out123_im),  
                             .Out124_re(Out124_re),  
                             .Out124_im(Out124_im),  
                             .Out125_re(Out125_re),  
                             .Out125_im(Out125_im),  
                             .Out126_re(Out126_re),  
                             .Out126_im(Out126_im),  
                             .Out127_re(Out127_re),  
                             .Out127_im(Out127_im),  
                             .Out128_re(Out128_re),  
                             .Out128_im(Out128_im)) ;
                                          initial begin
                                          clk=0;
                                          res=0;
                                          end
                                          always begin #5 clk=~clk; end
                                         
 initial begin                                         # 10 res=1;
 #20
                                        In128=11'b00011_000000;
  In129=11'b00011_000000;
  In130=11'b11101_000000;
  In131=11'b11101_000000;
  In132=11'b11011_000000;
  In133=11'b11011_000000;
  In134=11'b00101_000000;
  In135=11'b00101_000000;
  In136=11'b00101_101010;
  In137=11'b00101_101010;
  In138=11'b11010_010110;
  In139=11'b11010_010110;
  In140=11'b00001_011011;
  In141=11'b00001_011011;
  In142=11'b11110_100101;
  In143=11'b11110_100101;
  In144=11'b11000_100111;
  In145=11'b11000_100111;
  In146=11'b00111_011001;
  In147=11'b00111_011001;
  In148=11'b00011_000100;
  In149=11'b00011_000100;
  In150=11'b11100_111100;
  In151=11'b11100_111100;
  In152=11'b00000_110001;
  In153=11'b00000_110001;
  In154=11'b11111_001111;
  In155=11'b11111_001111;
  In156=11'b11110_001010;
  In157=11'b11110_001010;
  In158=11'b00001_110110;
  In159=11'b00001_110110;
  In160=11'b00100_110000;
  In161=11'b00100_110000;
  In162=11'b11011_010000;
  In163=11'b11011_010000;
  In164=11'b00101_101110;
  In165=11'b00101_101110;
  In166=11'b11010_010010;
  In167=11'b11010_010010;
  In168=11'b11101_100110;
  In169=11'b11101_100110;
  In170=11'b00010_011010;
  In171=11'b00010_011010;
  In172=11'b00010_101001;
  In173=11'b00010_101001;
  In174=11'b11101_010111;
  In175=11'b11101_010111;
  In176=11'b11111_010100;
  In177=11'b11111_010100;
  In178=11'b00000_101100;
  In179=11'b00000_101100;
  In180=11'b11000_100111;
  In181=11'b11000_100111;
  In182=11'b00111_011001;
  In183=11'b00111_011001;
  In184=11'b11111_110101;
  In185=11'b11111_110101;
  In186=11'b00000_001011;
  In187=11'b00000_001011;
  In188=11'b00011_100101;
  In189=11'b00011_100101;
  In190=11'b11100_011011;
  In191=11'b11100_011011;
  In192=11'b00110_101111;
  In193=11'b00110_101111;
  In194=11'b11001_010001;
  In195=11'b11001_010001;
  In196=11'b11111_100011;
  In197=11'b11111_100011;
  In198=11'b00000_011101;
  In199=11'b00000_011101;
  In200=11'b00001_100010;
  In201=11'b00001_100010;
  In202=11'b11110_011110;
  In203=11'b11110_011110;
  In204=11'b00100_011111;
  In205=11'b00100_011111;
  In206=11'b11011_100001;
  In207=11'b11011_100001;
  In208=11'b11001_010001;
  In209=11'b11001_010001;
  In210=11'b00110_101111;
  In211=11'b00110_101111;
  In212=11'b11011_111101;
  In213=11'b11011_111101;
  In214=11'b00100_000011;
  In215=11'b00100_000011;
  In216=11'b00010_010101;
  In217=11'b00010_010101;
  In218=11'b11101_101011;
  In219=11'b11101_101011;
  In220=11'b00000_111011;
  In221=11'b00000_111011;
  In222=11'b11111_000101;
  In223=11'b11111_000101;
  In224=11'b11110_000110;
  In225=11'b11110_000110;
  In226=11'b00001_111010;
  In227=11'b00001_111010;
  In228=11'b00111_101000;
  In229=11'b00111_101000;
  In230=11'b11000_011000;
  In231=11'b11000_011000;
  In232=11'b11101_101101;
  In233=11'b11101_101101;
  In234=11'b00010_010011;
  In235=11'b00010_010011;
  In236=11'b11111_000000;
  In237=11'b11111_000000;
  In238=11'b00001_000000;
  In239=11'b00001_000000;
  In240=11'b00101_000101;
  In241=11'b00101_000101;
  In242=11'b11010_111011;
  In243=11'b11010_111011;
  In244=11'b11011_100100;
  In245=11'b11011_100100;
  In246=11'b00100_011100;
  In247=11'b00100_011100;
  In248=11'b11011_101111;
  In249=11'b11011_101111;
  In250=11'b00100_010001;
  In251=11'b00100_010001;
  In252=11'b00010_000110;
  In253=11'b00010_000110;
  In254=11'b11101_111010;
  In255=11'b11101_111010;
                 
  #100;
  In128=11'b00000000000;
  In129=11'b00000000000;
  In130=11'b00000000000;
  In131=11'b00000000000;
  In132=11'b00000000000;
  In133=11'b00000000000;
  In134=11'b00000000000;
  In135=11'b00000000000;
  In136=11'b10000000000;
  In137=11'b10000000000;
  In138=11'b10000000000;
  In139=11'b10000000000;
  In140=11'b01111111111;
  In141=11'b01111111111;
  In142=11'b01111111111;
  In143=11'b01111111111;
  In144=11'b10100101100;
  In145=11'b10100101100;
  In146=11'b10100101100;
  In147=11'b10100101100;
  In148=11'b01011010100;
  In149=11'b01011010100;
  In150=11'b01011010100;
  In151=11'b01011010100;
  In152=11'b10100101100;
  In153=11'b10100101100;
  In154=11'b10100101100;
  In155=11'b10100101100;
  In156=11'b01011010100;
  In157=11'b01011010100;
  In158=11'b01011010100;
  In159=11'b01011010100;
  In160=11'b11001111000;
  In161=11'b11001111000;
  In162=11'b11001111000;
  In163=11'b11001111000;
  In164=11'b00110001000;
  In165=11'b00110001000;
  In166=11'b00110001000;
  In167=11'b00110001000;
  In168=11'b10001001110;
  In169=11'b10001001110;
  In170=11'b10001001110;
  In171=11'b10001001110;
  In172=11'b01110110010;
  In173=11'b01110110010;
  In174=11'b01110110010;
  In175=11'b01110110010;
  In176=11'b10001001110;
  In177=11'b10001001110;
  In178=11'b10001001110;
  In179=11'b10001001110;
  In180=11'b01110110010;
  In181=11'b01110110010;
  In182=11'b01110110010;
  In183=11'b01110110010;
  In184=11'b11001111000;
  In185=11'b11001111000;
  In186=11'b11001111000;
  In187=11'b11001111000;
  In188=11'b00110001000;
  In189=11'b00110001000;
  In190=11'b00110001000;
  In191=11'b00110001000;
  In192=11'b11100111000;
  In193=11'b11100111000;
  In194=11'b11100111000;
  In195=11'b11100111000;
  In196=11'b00011001000;
  In197=11'b00011001000;
  In198=11'b00011001000;
  In199=11'b00011001000;
  In200=11'b10000010100;
  In201=11'b10000010100;
  In202=11'b10000010100;
  In203=11'b10000010100;
  In204=11'b01111101100;
  In205=11'b01111101100;
  In206=11'b01111101100;
  In207=11'b01111101100;
  In208=11'b10010101101;
  In209=11'b10010101101;
  In210=11'b10010101101;
  In211=11'b10010101101;
  In212=11'b01101010011;
  In213=11'b01101010011;
  In214=11'b01101010011;
  In215=11'b01101010011;
  In216=11'b10111000111;
  In217=11'b10111000111;
  In218=11'b10111000111;
  In219=11'b10111000111;
  In220=11'b01000111001;
  In221=11'b01000111001;
  In222=11'b01000111001;
  In223=11'b01000111001;
  In224=11'b10111000111;
  In225=11'b10111000111;
  In226=11'b10111000111;
  In227=11'b10111000111;
  In228=11'b01000111001;
  In229=11'b01000111001;
  In230=11'b01000111001;
  In231=11'b01000111001;
  In232=11'b10010101101;
  In233=11'b10010101101;
  In234=11'b10010101101;
  In235=11'b10010101101;
  In236=11'b01101010011;
  In237=11'b01101010011;
  In238=11'b01101010011;
  In239=11'b01101010011;
  In240=11'b10000010100;
  In241=11'b10000010100;
  In242=11'b10000010100;
  In243=11'b10000010100;
  In244=11'b01111101100;
  In245=11'b01111101100;
  In246=11'b01111101100;
  In247=11'b01111101100;
  In248=11'b11100111000;
  In249=11'b11100111000;
  In250=11'b11100111000;
  In251=11'b11100111000;
  In252=11'b00011001000;
  In253=11'b00011001000;
  In254=11'b00011001000;
  In255=11'b00011001000;
  #100;
  In128=11'b11111111011;
  In129=11'b11111111011;
  In130=11'b11111111011;
  In131=11'b11111111011;
  In132=11'b00000000000;
  In133=11'b00000000000;
  In134=11'b00000000000;
  In135=11'b00000000000;
  In136=11'b00000000011;
  In137=11'b00000000011;
  In138=11'b00000000011;
  In139=11'b00000000011;
  In140=11'b11111111101;
  In141=11'b11111111101;
  In142=11'b11111111101;
  In143=11'b11111111101;
  In144=11'b11111111111;
  In145=11'b11111111111;
  In146=11'b11111111111;
  In147=11'b11111111111;
  In148=11'b00000000100;
  In149=11'b00000000100;
  In150=11'b00000000100;
  In151=11'b00000000100;
  In152=11'b11111111100;
  In153=11'b11111111100;
  In154=11'b11111111100;
  In155=11'b11111111100;
  In156=11'b00000000001;
  In157=11'b00000000001;
  In158=11'b00000000001;
  In159=11'b00000000001;
  In160=11'b11111111101;
  In161=11'b11111111101;
  In162=11'b11111111101;
  In163=11'b11111111101;
  In164=11'b00000000010;
  In165=11'b00000000010;
  In166=11'b00000000010;
  In167=11'b00000000010;
  In168=11'b00000000100;
  In169=11'b00000000100;
  In170=11'b00000000100;
  In171=11'b00000000100;
  In172=11'b11111111111;
  In173=11'b11111111111;
  In174=11'b11111111111;
  In175=11'b11111111111;
  In176=11'b00000000001;
  In177=11'b00000000001;
  In178=11'b00000000001;
  In179=11'b00000000001;
  In180=11'b11111111100;
  In181=11'b11111111100;
  In182=11'b11111111100;
  In183=11'b11111111100;
  In184=11'b11111111110;
  In185=11'b11111111110;
  In186=11'b11111111110;
  In187=11'b11111111110;
  In188=11'b00000000011;
  In189=11'b00000000011;
  In190=11'b00000000011;
  In191=11'b00000000011;
  In192=11'b11111111100;
  In193=11'b11111111100;
  In194=11'b11111111100;
  In195=11'b11111111100;
  In196=11'b00000000001;
  In197=11'b00000000001;
  In198=11'b00000000001;
  In199=11'b00000000001;
  In200=11'b00000000100;
  In201=11'b00000000100;
  In202=11'b00000000100;
  In203=11'b00000000100;
  In204=11'b11111111110;
  In205=11'b11111111110;
  In206=11'b11111111110;
  In207=11'b11111111110;
  In208=11'b00000000000;
  In209=11'b00000000000;
  In210=11'b00000000000;
  In211=11'b00000000000;
  In212=11'b00000000101;
  In213=11'b00000000101;
  In214=11'b00000000101;
  In215=11'b00000000101;
  In216=11'b11111111101;
  In217=11'b11111111101;
  In218=11'b11111111101;
  In219=11'b11111111101;
  In220=11'b00000000010;
  In221=11'b00000000010;
  In222=11'b00000000010;
  In223=11'b00000000010;
  In224=11'b11111111110;
  In225=11'b11111111110;
  In226=11'b11111111110;
  In227=11'b11111111110;
  In228=11'b00000000011;
  In229=11'b00000000011;
  In230=11'b00000000011;
  In231=11'b00000000011;
  In232=11'b11111111011;
  In233=11'b11111111011;
  In234=11'b11111111011;
  In235=11'b11111111011;
  In236=11'b00000000000;
  In237=11'b00000000000;
  In238=11'b00000000000;
  In239=11'b00000000000;
  In240=11'b00000000010;
  In241=11'b00000000010;
  In242=11'b00000000010;
  In243=11'b00000000010;
  In244=11'b11111111100;
  In245=11'b11111111100;
  In246=11'b11111111100;
  In247=11'b11111111100;
  In248=11'b11111111111;
  In249=11'b11111111111;
  In250=11'b11111111111;
  In251=11'b11111111111;
  In252=11'b00000000100;
  In253=11'b00000000100;
  In254=11'b00000000100;
  In255=11'b00000000100;
  #100;
  In128=11'b00000000000;
  In129=11'b00000000000;
  In130=11'b00000000000;
  In131=11'b00000000000;
  In132=11'b00000000000;
  In133=11'b00000000000;
  In134=11'b00000000000;
  In135=11'b00000000000;
  In136=11'b00111110010;
  In137=11'b00111110010;
  In138=11'b11000001110;
  In139=11'b11000001110;
  In140=11'b00000000000;
  In141=11'b00000000000;
  In142=11'b00000000000;
  In143=11'b00000000000;
  In144=11'b10101110110;
  In145=11'b10101110110;
  In146=11'b01010001010;
  In147=11'b01010001010;
  In148=11'b00000000000;
  In149=11'b00000000000;
  In150=11'b00000000000;
  In151=11'b00000000000;
  In152=11'b00100001101;
  In153=11'b00100001101;
  In154=11'b11011110011;
  In155=11'b11011110011;
  In156=11'b00000000000;
  In157=11'b00000000000;
  In158=11'b00000000000;
  In159=11'b00000000000;
  In160=11'b01001001001;
  In161=11'b01001001001;
  In162=11'b10110110111;
  In163=11'b10110110111;
  In164=11'b00000000000;
  In165=11'b00000000000;
  In166=11'b00000000000;
  In167=11'b00000000000;
  In168=11'b10101001110;
  In169=11'b10101001110;
  In170=11'b01010110010;
  In171=11'b01010110010;
  In172=11'b00000000000;
  In173=11'b00000000000;
  In174=11'b00000000000;
  In175=11'b00000000000;
  In176=11'b00010001001;
  In177=11'b00010001001;
  In178=11'b11101110111;
  In179=11'b11101110111;
  In180=11'b00000000000;
  In181=11'b00000000000;
  In182=11'b00000000000;
  In183=11'b00000000000;
  In184=11'b00110000111;
  In185=11'b00110000111;
  In186=11'b11001111001;
  In187=11'b11001111001;
  In188=11'b00000000000;
  In189=11'b00000000000;
  In190=11'b00000000000;
  In191=11'b00000000000;
  In192=11'b01001101101;
  In193=11'b01001101101;
  In194=11'b10110010011;
  In195=11'b10110010011;
  In196=11'b00000000000;
  In197=11'b00000000000;
  In198=11'b00000000000;
  In199=11'b00000000000;
  In200=11'b11100110100;
  In201=11'b11100110100;
  In202=11'b00011001100;
  In203=11'b00011001100;
  In204=11'b00000000000;
  In205=11'b00000000000;
  In206=11'b00000000000;
  In207=11'b00000000000;
  In208=11'b10111100000;
  In209=11'b10111100000;
  In210=11'b01000100000;
  In211=11'b01000100000;
  In212=11'b00000000000;
  In213=11'b00000000000;
  In214=11'b00000000000;
  In215=11'b00000000000;
  In216=11'b01010111101;
  In217=11'b01010111101;
  In218=11'b10101000011;
  In219=11'b10101000011;
  In220=11'b00000000000;
  In221=11'b00000000000;
  In222=11'b00000000000;
  In223=11'b00000000000;
  In224=11'b11110111011;
  In225=11'b11110111011;
  In226=11'b00001000101;
  In227=11'b00001000101;
  In228=11'b00000000000;
  In229=11'b00000000000;
  In230=11'b00000000000;
  In231=11'b00000000000;
  In232=11'b11001000001;
  In233=11'b11001000001;
  In234=11'b00110111111;
  In235=11'b00110111111;
  In236=11'b00000000000;
  In237=11'b00000000000;
  In238=11'b00000000000;
  In239=11'b00000000000;
  In240=11'b01010100010;
  In241=11'b01010100010;
  In242=11'b10101011110;
  In243=11'b10101011110;
  In244=11'b00000000000;
  In245=11'b00000000000;
  In246=11'b00000000000;
  In247=11'b00000000000;
  In248=11'b11010110100;
  In249=11'b11010110100;
  In250=11'b00101001100;
  In251=11'b00101001100;
  In252=11'b00000000000;
  In253=11'b00000000000;
  In254=11'b00000000000;
  In255=11'b00000000000;
  #100;
  In128=11'b00000000000;
  In129=11'b00000000000;
  In130=11'b00000000000;
  In131=11'b00000000000;
  In132=11'b00101011100;
  In133=11'b00101011100;
  In134=11'b11010100100;
  In135=11'b11010100100;
  In136=11'b11010101010;
  In137=11'b11010101010;
  In138=11'b11110101110;
  In139=11'b11110101110;
  In140=11'b00001010010;
  In141=11'b00001010010;
  In142=11'b00101010110;
  In143=11'b00101010110;
  In144=11'b00101100000;
  In145=11'b00101100000;
  In146=11'b11100000010;
  In147=11'b11100000010;
  In148=11'b11100001111;
  In149=11'b11100001111;
  In150=11'b11010100000;
  In151=11'b11010100000;
  In152=11'b00101100000;
  In153=11'b00101100000;
  In154=11'b00011110001;
  In155=11'b00011110001;
  In156=11'b00011111110;
  In157=11'b00011111110;
  In158=11'b11010100000;
  In159=11'b11010100000;
  In160=11'b11010100001;
  In161=11'b11010100001;
  In162=11'b00001110100;
  In163=11'b00001110100;
  In164=11'b00100010001;
  In165=11'b00100010001;
  In166=11'b00100110110;
  In167=11'b00100110110;
  In168=11'b00101100000;
  In169=11'b00101100000;
  In170=11'b11010111011;
  In171=11'b11010111011;
  In172=11'b11101111011;
  In173=11'b11101111011;
  In174=11'b11100001000;
  In175=11'b11100001000;
  In176=11'b00011111000;
  In177=11'b00011111000;
  In178=11'b00010000101;
  In179=11'b00010000101;
  In180=11'b00101000101;
  In181=11'b00101000101;
  In182=11'b11010100000;
  In183=11'b11010100000;
  In184=11'b11011001010;
  In185=11'b11011001010;
  In186=11'b11011101111;
  In187=11'b11011101111;
  In188=11'b11110001100;
  In189=11'b11110001100;
  In190=11'b00101011111;
  In191=11'b00101011111;
  In192=11'b11100111110;
  In193=11'b11100111110;
  In194=11'b00101100000;
  In195=11'b00101100000;
  In196=11'b11010110011;
  In197=11'b11010110011;
  In198=11'b11011100111;
  In199=11'b11011100111;
  In200=11'b00011000000;
  In201=11'b00011000000;
  In202=11'b00101000011;
  In203=11'b00101000011;
  In204=11'b11010100000;
  In205=11'b11010100000;
  In206=11'b00100101001;
  In207=11'b00100101001;
  In208=11'b00000010101;
  In209=11'b00000010101;
  In210=11'b11010100011;
  In211=11'b11010100011;
  In212=11'b00101001010;
  In213=11'b00101001010;
  In214=11'b00010111000;
  In215=11'b00010111000;
  In216=11'b11010101011;
  In217=11'b11010101011;
  In218=11'b00101011111;
  In219=11'b00101011111;
  In220=11'b11101111001;
  In221=11'b11101111001;
  In222=11'b11110111011;
  In223=11'b11110111011;
  In224=11'b00001000101;
  In225=11'b00001000101;
  In226=11'b00010000111;
  In227=11'b00010000111;
  In228=11'b11010100001;
  In229=11'b11010100001;
  In230=11'b00101010101;
  In231=11'b00101010101;
  In232=11'b11101001000;
  In233=11'b11101001000;
  In234=11'b11010110110;
  In235=11'b11010110110;
  In236=11'b00101011101;
  In237=11'b00101011101;
  In238=11'b11111101011;
  In239=11'b11111101011;
  In240=11'b11011010111;
  In241=11'b11011010111;
  In242=11'b00101100000;
  In243=11'b00101100000;
  In244=11'b11010111101;
  In245=11'b11010111101;
  In246=11'b11101000000;
  In247=11'b11101000000;
  In248=11'b00100011001;
  In249=11'b00100011001;
  In250=11'b00101001101;
  In251=11'b00101001101;
  In252=11'b11010100000;
  In253=11'b11010100000;
  In254=11'b00011000010;
  In255=11'b00011000010;
#100  $finish;
  end                             
endmodule
